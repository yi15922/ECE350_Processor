module inverter(out, in); 
    input [31:0] in; 
    output [31:0] out; 

    not invert0(out[0], in[0]); 
    not invert1(out[1], in[1]); 
    not invert2(out[2], in[2]); 
    not invert3(out[3], in[3]); 
    not invert4(out[4], in[4]); 
    not invert5(out[5], in[5]); 
    not invert6(out[6], in[6]); 
    not invert7(out[7], in[7]); 
    not invert8(out[8], in[8]); 
    not invert9(out[9], in[9]); 
    not invert10(out[10], in[10]); 
    not invert11(out[11], in[11]); 
    not invert12(out[12], in[12]); 
    not invert13(out[13], in[13]); 
    not invert14(out[14], in[14]); 
    not invert15(out[15], in[15]); 
    not invert16(out[16], in[16]); 
    not invert17(out[17], in[17]); 
    not invert18(out[18], in[18]); 
    not invert19(out[19], in[19]); 
    not invert20(out[20], in[20]); 
    not invert21(out[21], in[21]); 
    not invert22(out[22], in[22]); 
    not invert23(out[23], in[23]); 
    not invert24(out[24], in[24]); 
    not invert25(out[25], in[25]); 
    not invert26(out[26], in[26]); 
    not invert27(out[27], in[27]); 
    not invert28(out[28], in[28]); 
    not invert29(out[29], in[29]); 
    not invert30(out[30], in[30]); 
    not invert31(out[31], in[31]); 


endmodule